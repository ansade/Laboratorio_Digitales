`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:30:52 01/30/2011
// Design Name:   MiniAlu
// Module Name:   D:/Proyecto/RTL/Dev/MiniALU/TestBench.v
// Project Name:  MiniALU
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: MiniAlu
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TestBench;

	// Inputs
	reg Clock;
	reg Reset;
	reg Reset2;

	// Outputs
	wire [7:0] oLed;

	// Instantiate the Unit Under Test (UUT)
	MiniAlu uut (
		.Clock(Clock), 
		.Reset(Reset), 
		.oLed(oLed),
		.Reset2(Reset2)
	);
	
	always
	begin
		#5  Clock =  ! Clock;
	end

	initial begin
		// Initialize Inputs
		Clock  = 0;
		Reset  = 0;
		Reset2 = 0;

		// Wait 100 ns for global reset to finish
		#50
		Reset2 = 1;
		#50
		Reset2 = 0;		
		#50;
		Reset = 1;
		#100
		Reset = 0;
        
		// Add stimulus here

	end
      
endmodule

